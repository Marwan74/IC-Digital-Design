module UART_wrapper (clk, rst, din, tx_wr_en, rx_rd_en, rx, dout, tx, framing_error, rx_empty, rx_full, tx_full);
    parameter WIDTH = 8;

    input clk, rst;
    input rx_rd_en; // Read enable for RX FIFO
    input tx_wr_en; // WRITE enable for TX FIFO
    input rx;       // Serial in
    input [WIDTH - 1 : 0] din; // Data to Transmit

    output rx_empty,rx_full; // RX FIFO status
    output tx_full;          // TX FIFO status
    output [WIDTH - 1 : 0] dout; // Data read from RX FIFO
    output tx;               // Serial out
    output framing_error;    // Error flag from RX

    // --- Internal Wires ---
    // These wires connect the sub-modules together.
   wire S_tick;         // The sample tick generated by the Baud_Generator

    // Baud rate generator
    Baud_Generator baud (.clk(clk), .rst(rst), .sample_tick(S_tick));

    // Tranmitter Top
    Transmitter_TOP tx_top (.clk(clk), .rst(rst), .S_tick(S_tick), .tx_wr_data(din), .tx_wr_en(tx_wr_en),
                           .tx(tx), .tx_full(tx_full));

    // Receiver Top
    Receiver_TOP rx_top (.clk(clk), .rst(rst), .S_tick(S_tick), .rx(rx), .rx_rd_en(rx_rd_en), .rx_rd_data(dout),
                         .rx_empty(rx_empty), .rx_full(rx_full), .frame_error(framing_error));
endmodule
